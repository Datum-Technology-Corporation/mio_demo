// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_CONSTANTS_SV__
`define __UVME_MAPU_CONSTANTS_SV__


const int unsigned  uvme_mapu_default_num_items_cons = 10; ///< Default number of Sequence Items to be generated in a Sequence.


`endif // __UVME_MAPU_CONSTANTS_SV__