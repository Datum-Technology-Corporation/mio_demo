// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_DADDER_DP_OUT_IF_CHKR_SV__
`define __UVMA_DADDER_DP_OUT_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_dadder_dp_out_if.
 * This module must be bound to an interface in a test bench.
 * @ingroup uvma_dadder_dp_out_misc
 */
module uvma_dadder_dp_out_if_chkr (
   uvma_dadder_dp_out_if  dadder_dp_out_if
);

   // TODO Add assertions to uvma_dadder_dp_out_if_chkr

endmodule : uvma_dadder_dp_out_if_chkr


`endif // __UVMA_DADDER_DP_OUT_IF_CHKR_SV__