// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __MAPU_MACROS_SVH__
`define __MAPU_MACROS_SVH__


`define MAPU_OP_ADD  2'b00
`define MAPU_OP_MULT 2'b01


`endif // __MAPU_MACROS_SVH__
