// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_MACROS_SVH__
`define __UVMA_MAPU_MACROS_SVH__


`ifndef UVMA_MAPU_MAX_DATA_WIDTH
   `define UVMA_MAPU_MAX_DATA_WIDTH 64
`endif


`endif // __UVMA_MAPU_MACROS_SVH__
