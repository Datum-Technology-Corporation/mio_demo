// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_DADDER_DP_OUT_TDEFS_SV__
`define __UVMA_DADDER_DP_OUT_TDEFS_SV__


typedef bit   [(`UVMA_DADDER_DP_OUT_MAX_DATA_WIDTH-1):0]  uvma_dadder_dp_out_data_b_t;
typedef logic [(`UVMA_DADDER_DP_OUT_MAX_DATA_WIDTH-1):0]  uvma_dadder_dp_out_data_l_t;


`endif // __UVMA_DADDER_DP_OUT_TDEFS_SV__