// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_DADDER_CONSTANTS_SV__
`define __UVME_DADDER_CONSTANTS_SV__


const int unsigned  uvme_dadder_default_clk_frequency = 100_000_000; ///< Clock agent frequency (Hz)
const int unsigned  uvme_dadder_default_data_width    =           8; ///< Data bus width in bits (b)


`endif // __UVME_DADDER_CONSTANTS_SV__