// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_DADDER_DP_IN_CONSTANTS_SV__
`define __UVMA_DADDER_DP_IN_CONSTANTS_SV__


const int unsigned  uvma_dadder_dp_in_default_data_width = 8;


`endif // __UVMA_DADDER_DP_IN_CONSTANTS_SV__