// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_IF_CHKR_SV__
`define __UVMA_MAPU_IF_CHKR_SV__


/**
 * Module encapsulating assertions targeting Matrix APU Block Agent interface.
 * @ingroup uvma_mapu_misc
 */
module uvma_mapu_if_chkr (
   uvma_mapu_if  agent_if ///< Target interface
);

   // TODO Add assertions to uvme_mapu_chkr

endmodule : uvma_mapu_if_chkr


`endif // __UVMA_MAPU_IF_CHKR_SV__