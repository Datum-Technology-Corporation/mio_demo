// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_DADDER_CP_TDEFS_SV__
`define __UVMA_DADDER_CP_TDEFS_SV__


/**
 * Valid operations.
 */
typedef enum bit {
   UVMA_DADDER_CP_OP_ADD      = 1,
   UVMA_DADDER_CP_OP_SUBTRACT = 0
} uvma_dadder_cp_op_enum;


`endif // __UVMA_DADDER_CP_TDEFS_SV__