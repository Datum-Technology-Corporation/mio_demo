// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_DADDER_MACROS_SVH__
`define __UVMT_DADDER_MACROS_SVH__


`ifndef UVMT_DADDER_DATA_WIDTH
   `define UVMT_DADDER_DATA_WIDTH 8
`endif


`endif // __UVMT_DADDER_MACROS_SVH__