// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __MAPU_MACROS_SVH__
`define __MAPU_MACROS_SVH__


`define MAPU_OP_ADD  1'b0
`define MAPU_OP_MULT 1'b1


`endif // __MAPU_MACROS_SVH__
