// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_MACROS_SVH__
`define __UVME_MAPU_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_MAPU_ABC
//        `define UVME_MAPU_ABC 32
//     `endif


`endif // __UVME_MAPU_MACROS_SVH__