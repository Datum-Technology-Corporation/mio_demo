// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_DADDER_TDEFS_SV__
`define __UVMT_DADDER_TDEFS_SV__


// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVMT_DADDER_ABC_MAX_WIDTH-1):0]  uvmt_dadder_abc_b_t;
// Ex: typedef enum {
//        UVMT_DADDER_MY_ABC
//     } uvmt_dadder_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_dadder_my_struct;


`endif // __UVMT_DADDER_TDEFS_SV__