// Copyright 2022 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_CONSTANTS_SV__
`define __UVMA_MAPU_CONSTANTS_SV__


const int unsigned  uvma_mapu_default_data_width = 32;


`endif // __UVMA_MAPU_CONSTANTS_SV__
