// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_MACROS_SVH__
`define __UVMT_MAPU_MACROS_SVH__


`ifndef UVMT_MAPU_DATA_WIDTH
   `define UVMT_MAPU_DATA_WIDTH 32
`endif


`endif // __UVMT_MAPU_MACROS_SVH__