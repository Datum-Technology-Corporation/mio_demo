// Copyright 2022 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_CONSTANTS_SV__
`define __UVMA_MAPU_CONSTANTS_SV__


// Add constants here
// Ex: const int unsigned  uvma_mapu_my_cons = 10;


`endif // __UVMA_MAPU_CONSTANTS_SV__