// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_DADDER_CP_MACROS_SVH__
`define __UVMA_DADDER_CP_MACROS_SVH__


`ifndef UVMA_DADDER_CP_MAX_DATA_WIDTH
   `define UVMA_DADDER_CP_MAX_DATA_WIDTH 32
`endif


`endif // __UVMA_DADDER_CP_MACROS_SVH__