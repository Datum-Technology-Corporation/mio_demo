// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_MACROS_SVH__
`define __UVMT_MAPU_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_MAPU_ABC_MAX_WIDTH
//        `define UVMT_MAPU_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMT_MAPU_MACROS_SVH__