// Copyright 2022 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_TDEFS_SV__
`define __UVMT_MAPU_TDEFS_SV__


// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVMT_MAPU_ABC_MAX_WIDTH-1):0]  uvmt_mapu_abc_b_t;
// Ex: typedef enum {
//        UVMT_MAPU_MY_ABC
//     } uvmt_mapu_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_mapu_my_struct;


`endif // __UVMT_MAPU_TDEFS_SV__