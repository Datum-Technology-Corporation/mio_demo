// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MAPU_MACROS_SVH__
`define __UVMA_MAPU_MACROS_SVH__


`define UVMA_MAPU_DATA_MAX_WIDTH  32



`endif // __UVMA_MAPU_MACROS_SVH__