// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_DADDER_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_DADDER_BASE_TEST_WORKAROUNDS_SV__


// Temporary configuration constraints here (this file should be empty by the end of the project).


`endif // __UVMT_DADDER_BASE_TEST_WORKAROUNDS_SV__