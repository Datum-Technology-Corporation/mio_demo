// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __MAPU_TDEFS_SV__
`define __MAPU_TDEFS_SV__





`endif // __MAPU_TDEFS_SV__
