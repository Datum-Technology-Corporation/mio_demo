// Copyright 2023 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MAPU_CONSTANTS_SV__
`define __UVME_MAPU_CONSTANTS_SV__


// Add constants here
// Ex: const int unsigned  uvme_mapu_example_cons = 10;


`endif // __UVME_MAPU_CONSTANTS_SV__