// Copyright 2022 Contributors
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_DADDER_MACROS_SVH__
`define __UVME_DADDER_MACROS_SVH__


`ifndef UVME_DADDER_MAX_DATA_WIDTH
   `define UVME_DADDER_MAX_DATA_WIDTH 32
`endif


`endif // __UVME_DADDER_MACROS_SVH__