// Copyright 2022 Acme Enterprises Inc.
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_MAPU_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_MAPU_BASE_TEST_WORKAROUNDS_SV__


// Temporary configuration constraints here (this file should be empty by the end of the project).


`endif // __UVMT_MAPU_BASE_TEST_WORKAROUNDS_SV__